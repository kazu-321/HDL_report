// 分周器(100Hz)
module m_prescale(input clk,output c_out);
	reg [19:0] cnt;
	wire wcout;
	
	assign wcout=(cnt==20'd499999) ? 1'b1 : 1'b0;
	assign c_out=wcout;
	
	always @(posedge clk) begin
		if (wcout)
			cnt <= 20'd0;
		else
			cnt <= cnt + 20'd1;
	end

endmodule


module m_matrix_key(
	input             clk, rst,	// クロック，リセット
	input      [3:0]  row, 			// 4bit入力 行
	output reg [3:0]  col,			// 4bit出力 列
	output reg [15:0] key,			// 16bitキー出力
	output            tc				// 出力カウント
	) ;
	
	reg [2:0]  index ;	
	reg [15:0] tmp ;

	always @(posedge rst or posedge clk) begin
		if(rst == 1'b1)begin
		   tmp   <= 16'hFFFF ;
			key   <= 16'h0000 ;
			index <= 3'd0 ;
		end
		else begin
			//LSB=0 colへの出力をセット
			if (index[0] == 1'b0) begin
				case (index[2:1]) 
					2'd0: begin
								col <= 4'b1110 ;
								key <= ~tmp ;
								tmp <= 16'hFFFF ;
							end
					2'd1: col <= 4'b1101 ;
					2'd2: col <= 4'b1011 ;
					2'd3: col <= 4'b0111 ;
				endcase
			end
			//LSB=1 rowの値を読む
			else begin
				tmp[{2'd0, index[2:1]}] <= row[0] ;
				tmp[{2'd1, index[2:1]}] <= row[1] ;
				tmp[{2'd2, index[2:1]}] <= row[2] ;
				tmp[{2'd3, index[2:1]}] <= row[3] ;
			end
			
			index <= index + 3'd1 ;		
			
		end
	end
	
	assign tc = (index == 3'd0) ? 1'b1 : 1'b0 ;
	 
endmodule

// 16bit→4bitデコーダ(計算機仕様に変更)
module m_dec16to4_calc (
    input [15:0] key,		// 16bit入力
    output [3:0] out,		// 4bit出力
    output       pushed		//打鍵検出
) ;

    function [4:0] f ;
        input [15:0] in ;
        case(in)
			  16'h0001: f = { 1'b1, 4'h1 } ;		// 0000_0000_0000_0001 → 4'h1
			  16'h0002: f = { 1'b1, 4'h2 } ;		// 0000_0000_0000_0010 → 4'h2
			  16'h0004: f = { 1'b1, 4'h3 } ;		// 0000_0000_0000_0100 → 4'h3
			  16'h0008: f = { 1'b1, 4'hA } ;		// 0000_0000_0000_1000 → 4'hA
			  16'h0010: f = { 1'b1, 4'h4 } ;		// 0000_0000_0001_0000 → 4'h4
			  16'h0020: f = { 1'b1, 4'h5 } ;		// 0000_0000_0010_0000 → 4'h5
			  16'h0040: f = { 1'b1, 4'h6 } ;		// 0000_0000_0100_0000 → 4'h6
			  16'h0080: f = { 1'b1, 4'hB } ;		// 0000_0000_1000_0000 → 4'hB
			  16'h0100: f = { 1'b1, 4'h7 } ;		// 0000_0001_0000_0000 → 4'h7
			  16'h0200: f = { 1'b1, 4'h8 } ;		// 0000_0010_0000_0000 → 4'h8
			  16'h0400: f = { 1'b1, 4'h9 } ;		// 0000_0100_0000_0000 → 4'h9
			  16'h0800: f = { 1'b1, 4'hC } ;		// 0000_1000_0000_0000 → 4'hC
			  16'h1000: f = { 1'b1, 4'hE } ;		// 0001_0000_0000_0000 → 4'hE
			  16'h2000: f = { 1'b1, 4'h0 } ;		// 0010_0000_0000_0000 → 4'h0
			  16'h4000: f = { 1'b1, 4'hF } ;		// 0100_0000_0000_0000 → 4'hF
			  16'h8000: f = { 1'b1, 4'hD } ;		// 1000_0000_0000_0000 → 4'hD
			  default:  f = { 1'b0, 4'h0 } ;		// キーが一つだけ押されているとき以外は pushed=0, out=0
        endcase
    endfunction

    assign { pushed, out } = f(key) ;

endmodule

